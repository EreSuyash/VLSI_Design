magic
tech sky130A
timestamp 1726439019
<< nwell >>
rect -31 127 0 284
rect 307 127 969 283
rect -65 -214 23 -61
rect -84 -218 23 -214
rect 176 -218 232 -61
rect 384 -218 445 -61
rect 577 -218 1045 -61
<< nmos >>
rect 748 47 763 89
rect 867 47 882 89
rect 770 -305 785 -263
rect 978 -305 993 -263
<< pmos >>
rect 748 147 763 265
rect 867 147 882 265
rect 770 -198 785 -80
rect 978 -198 993 -80
<< ndiff >>
rect 714 80 748 89
rect 714 63 720 80
rect 737 63 748 80
rect 714 47 748 63
rect 763 81 797 89
rect 763 64 772 81
rect 789 64 797 81
rect 763 47 797 64
rect 833 81 867 89
rect 833 64 841 81
rect 858 64 867 81
rect 833 47 867 64
rect 882 80 916 89
rect 882 63 893 80
rect 910 63 916 80
rect 882 47 916 63
rect 736 -272 770 -263
rect 736 -289 742 -272
rect 759 -289 770 -272
rect 736 -305 770 -289
rect 785 -271 819 -263
rect 785 -288 794 -271
rect 811 -288 819 -271
rect 785 -305 819 -288
rect 944 -272 978 -263
rect 944 -289 950 -272
rect 967 -289 978 -272
rect 944 -305 978 -289
rect 993 -271 1027 -263
rect 993 -288 1002 -271
rect 1019 -288 1027 -271
rect 993 -305 1027 -288
<< pdiff >>
rect 714 246 748 265
rect 714 229 721 246
rect 738 229 748 246
rect 714 212 748 229
rect 714 195 721 212
rect 738 195 748 212
rect 714 178 748 195
rect 714 161 720 178
rect 737 161 748 178
rect 714 147 748 161
rect 763 246 797 265
rect 763 229 773 246
rect 790 229 797 246
rect 763 212 797 229
rect 763 195 773 212
rect 790 195 797 212
rect 763 178 797 195
rect 763 161 773 178
rect 790 161 797 178
rect 763 147 797 161
rect 833 246 867 265
rect 833 229 840 246
rect 857 229 867 246
rect 833 212 867 229
rect 833 195 840 212
rect 857 195 867 212
rect 833 178 867 195
rect 833 161 840 178
rect 857 161 867 178
rect 833 147 867 161
rect 882 246 916 265
rect 882 229 892 246
rect 909 229 916 246
rect 882 212 916 229
rect 882 195 892 212
rect 909 195 916 212
rect 882 178 916 195
rect 882 161 893 178
rect 910 161 916 178
rect 882 147 916 161
rect 736 -99 770 -80
rect 736 -116 743 -99
rect 760 -116 770 -99
rect 736 -133 770 -116
rect 736 -150 743 -133
rect 760 -150 770 -133
rect 736 -167 770 -150
rect 736 -184 742 -167
rect 759 -184 770 -167
rect 736 -198 770 -184
rect 785 -99 819 -80
rect 785 -116 795 -99
rect 812 -116 819 -99
rect 785 -133 819 -116
rect 785 -150 795 -133
rect 812 -150 819 -133
rect 785 -167 819 -150
rect 785 -184 795 -167
rect 812 -184 819 -167
rect 785 -198 819 -184
rect 944 -99 978 -80
rect 944 -116 951 -99
rect 968 -116 978 -99
rect 944 -133 978 -116
rect 944 -150 951 -133
rect 968 -150 978 -133
rect 944 -167 978 -150
rect 944 -184 950 -167
rect 967 -184 978 -167
rect 944 -198 978 -184
rect 993 -99 1027 -80
rect 993 -116 1003 -99
rect 1020 -116 1027 -99
rect 993 -133 1027 -116
rect 993 -150 1003 -133
rect 1020 -150 1027 -133
rect 993 -167 1027 -150
rect 993 -184 1003 -167
rect 1020 -184 1027 -167
rect 993 -198 1027 -184
<< ndiffc >>
rect 720 63 737 80
rect 772 64 789 81
rect 841 64 858 81
rect 893 63 910 80
rect 742 -289 759 -272
rect 794 -288 811 -271
rect 950 -289 967 -272
rect 1002 -288 1019 -271
<< pdiffc >>
rect 721 229 738 246
rect 721 195 738 212
rect 720 161 737 178
rect 773 229 790 246
rect 773 195 790 212
rect 773 161 790 178
rect 840 229 857 246
rect 840 195 857 212
rect 840 161 857 178
rect 892 229 909 246
rect 892 195 909 212
rect 893 161 910 178
rect 743 -116 760 -99
rect 743 -150 760 -133
rect 742 -184 759 -167
rect 795 -116 812 -99
rect 795 -150 812 -133
rect 795 -184 812 -167
rect 951 -116 968 -99
rect 951 -150 968 -133
rect 950 -184 967 -167
rect 1003 -116 1020 -99
rect 1003 -150 1020 -133
rect 1003 -184 1020 -167
<< psubdiff >>
rect 699 -276 736 -263
rect 699 -293 708 -276
rect 725 -293 736 -276
rect 699 -305 736 -293
rect 907 -276 944 -263
rect 907 -293 916 -276
rect 933 -293 944 -276
rect 907 -305 944 -293
<< nsubdiff >>
rect 702 -127 736 -80
rect 702 -144 709 -127
rect 726 -144 736 -127
rect 702 -198 736 -144
rect 910 -127 944 -80
rect 910 -144 917 -127
rect 934 -144 944 -127
rect 910 -198 944 -144
<< psubdiffcont >>
rect 708 -293 725 -276
rect 916 -293 933 -276
<< nsubdiffcont >>
rect 709 -144 726 -127
rect 917 -144 934 -127
<< poly >>
rect 87 299 882 317
rect 87 278 102 299
rect 748 265 763 278
rect 867 265 882 299
rect 748 139 763 147
rect 147 123 206 138
rect 664 132 763 139
rect 867 139 882 147
rect 867 138 966 139
rect 21 -17 36 107
rect 147 28 162 123
rect 305 107 406 122
rect 664 115 672 132
rect 689 123 763 132
rect 808 131 966 138
rect 808 123 941 131
rect 689 115 697 123
rect 664 107 697 115
rect 111 13 162 28
rect -13 -22 36 -17
rect 197 -22 212 0
rect -13 -37 212 -22
rect -13 -214 3 -37
rect -83 -222 4 -214
rect -224 -247 -165 -232
rect -83 -239 -75 -222
rect -58 -229 4 -222
rect -58 -239 -50 -229
rect -83 -247 -50 -239
rect -224 -340 -209 -247
rect 391 -340 406 107
rect 682 -17 697 107
rect 748 89 763 102
rect 748 28 763 47
rect 808 28 823 123
rect 933 114 941 123
rect 958 114 966 131
rect 933 107 966 114
rect 867 89 882 102
rect 867 28 882 47
rect 739 23 823 28
rect 739 6 747 23
rect 764 13 823 23
rect 852 19 885 28
rect 764 6 772 13
rect 739 0 772 6
rect 852 2 860 19
rect 877 2 885 19
rect 648 -22 697 -17
rect 852 -5 885 2
rect 852 -22 873 -5
rect 648 -37 873 -22
rect 648 -214 664 -37
rect 770 -80 785 -67
rect 978 -80 993 -67
rect 770 -214 785 -198
rect 978 -214 993 -198
rect 648 -340 665 -214
rect 737 -222 785 -214
rect 737 -239 745 -222
rect 762 -239 785 -222
rect 737 -247 785 -239
rect 945 -222 993 -214
rect 945 -239 953 -222
rect 970 -239 993 -222
rect 945 -247 993 -239
rect 770 -263 785 -247
rect 978 -263 993 -247
rect 770 -318 785 -305
rect 978 -318 993 -305
rect -224 -355 665 -340
<< polycont >>
rect 672 115 689 132
rect -75 -239 -58 -222
rect 941 114 958 131
rect 747 6 764 23
rect 860 2 877 19
rect 745 -239 762 -222
rect 953 -239 970 -222
<< locali >>
rect -220 277 -185 294
rect -220 -52 -203 277
rect 714 246 745 265
rect 714 229 721 246
rect 738 229 745 246
rect 714 212 745 229
rect 714 195 721 212
rect 738 195 745 212
rect 714 178 745 195
rect 714 161 720 178
rect 737 161 745 178
rect 664 132 697 139
rect -131 98 -130 131
rect 664 115 672 132
rect 689 115 697 132
rect 664 107 697 115
rect 714 80 745 161
rect 714 64 720 80
rect -48 47 54 64
rect 136 47 172 64
rect 255 47 418 64
rect 146 -17 163 47
rect -13 -34 163 -17
rect -166 -247 -165 -214
rect -83 -222 -50 -214
rect -83 -239 -75 -222
rect -58 -239 -50 -222
rect -83 -247 -50 -239
rect -13 -228 4 -34
rect 401 -87 418 47
rect 614 63 720 64
rect 737 63 745 80
rect 614 47 745 63
rect 766 246 797 258
rect 766 229 773 246
rect 790 229 797 246
rect 766 212 797 229
rect 766 195 773 212
rect 790 195 797 212
rect 766 178 797 195
rect 766 161 773 178
rect 790 161 797 178
rect 766 81 797 161
rect 766 64 772 81
rect 789 64 797 81
rect 833 246 864 258
rect 833 229 840 246
rect 857 229 864 246
rect 833 212 864 229
rect 833 195 840 212
rect 857 195 864 212
rect 833 178 864 195
rect 833 161 840 178
rect 857 161 864 178
rect 833 81 864 161
rect 833 64 841 81
rect 858 64 864 81
rect 766 47 864 64
rect 885 246 916 265
rect 885 229 892 246
rect 909 229 916 246
rect 885 212 916 229
rect 885 195 892 212
rect 909 195 916 212
rect 885 178 916 195
rect 885 161 893 178
rect 910 161 916 178
rect 885 80 916 161
rect 933 131 966 139
rect 933 114 941 131
rect 958 114 966 131
rect 933 107 966 114
rect 885 63 893 80
rect 910 64 916 80
rect 910 63 1079 64
rect 885 47 1079 63
rect 614 -87 631 47
rect 739 23 772 28
rect 739 6 747 23
rect 764 6 772 23
rect 739 0 772 6
rect 807 -17 824 47
rect 852 19 885 28
rect 852 2 860 19
rect 877 2 885 19
rect 852 -5 885 2
rect 366 -104 418 -87
rect 572 -104 631 -87
rect 648 -34 824 -17
rect -13 -245 76 -228
rect 158 -240 284 -223
rect 648 -228 665 -34
rect 682 -68 689 -51
rect 706 -68 770 -51
rect 787 -68 814 -51
rect 831 -68 837 -51
rect 890 -68 897 -51
rect 914 -68 978 -51
rect 995 -68 1022 -51
rect 1039 -68 1045 -51
rect 736 -85 767 -68
rect 944 -85 975 -68
rect 702 -99 767 -85
rect 702 -116 743 -99
rect 760 -116 767 -99
rect 702 -127 767 -116
rect 702 -144 709 -127
rect 726 -133 767 -127
rect 726 -144 743 -133
rect 702 -150 743 -144
rect 760 -150 767 -133
rect 702 -167 767 -150
rect 702 -184 742 -167
rect 759 -184 767 -167
rect 702 -192 767 -184
rect 788 -99 819 -87
rect 788 -116 795 -99
rect 812 -116 819 -99
rect 788 -133 819 -116
rect 788 -150 795 -133
rect 812 -150 819 -133
rect 788 -167 819 -150
rect 788 -184 795 -167
rect 812 -184 819 -167
rect 737 -222 770 -214
rect 737 -228 745 -222
rect 195 -356 212 -240
rect 401 -247 490 -230
rect 648 -239 745 -228
rect 762 -239 770 -222
rect 648 -245 770 -239
rect 737 -247 770 -245
rect 788 -223 819 -184
rect 910 -99 975 -85
rect 1062 -87 1079 47
rect 910 -116 951 -99
rect 968 -116 975 -99
rect 910 -127 975 -116
rect 910 -144 917 -127
rect 934 -133 975 -127
rect 934 -144 951 -133
rect 910 -150 951 -144
rect 968 -150 975 -133
rect 910 -167 975 -150
rect 910 -184 950 -167
rect 967 -184 975 -167
rect 910 -192 975 -184
rect 996 -99 1079 -87
rect 996 -116 1003 -99
rect 1020 -104 1079 -99
rect 1020 -116 1027 -104
rect 996 -133 1027 -116
rect 996 -150 1003 -133
rect 1020 -150 1027 -133
rect 996 -167 1027 -150
rect 996 -184 1003 -167
rect 1020 -184 1027 -167
rect 945 -222 978 -214
rect 945 -223 953 -222
rect 788 -239 953 -223
rect 970 -239 978 -222
rect 788 -240 978 -239
rect 401 -356 418 -247
rect 701 -272 767 -265
rect 701 -276 742 -272
rect 701 -293 708 -276
rect 725 -289 742 -276
rect 759 -289 767 -272
rect 725 -293 767 -289
rect 701 -305 767 -293
rect 788 -271 819 -240
rect 853 -241 870 -240
rect 945 -247 978 -240
rect 788 -288 794 -271
rect 811 -288 819 -271
rect 788 -305 819 -288
rect 909 -272 975 -265
rect 909 -276 950 -272
rect 909 -293 916 -276
rect 933 -289 950 -276
rect 967 -289 975 -272
rect 933 -293 975 -289
rect 909 -305 975 -293
rect 996 -271 1027 -184
rect 996 -288 1002 -271
rect 1019 -288 1027 -271
rect 996 -305 1027 -288
rect 736 -322 767 -305
rect 944 -322 975 -305
rect 682 -339 690 -322
rect 707 -339 770 -322
rect 787 -339 814 -322
rect 831 -339 837 -322
rect 890 -339 898 -322
rect 915 -339 978 -322
rect 995 -339 1022 -322
rect 1039 -339 1045 -322
rect 195 -373 418 -356
<< viali >>
rect 689 -68 706 -51
rect 770 -68 787 -51
rect 814 -68 831 -51
rect 897 -68 914 -51
rect 978 -68 995 -51
rect 1022 -68 1039 -51
rect 690 -339 707 -322
rect 770 -339 787 -322
rect 814 -339 831 -322
rect 898 -339 915 -322
rect 978 -339 995 -322
rect 1022 -339 1039 -322
<< metal1 >>
rect -186 274 -185 297
rect -292 3 -185 26
rect -292 -319 -262 3
rect -65 -71 21 -48
rect 176 -71 229 -48
rect 646 -49 1045 -48
rect 384 -51 1045 -49
rect 384 -68 689 -51
rect 706 -68 770 -51
rect 787 -68 814 -51
rect 831 -68 897 -51
rect 914 -68 978 -51
rect 995 -68 1022 -51
rect 1039 -68 1045 -51
rect 384 -71 1045 -68
rect -292 -342 -220 -319
rect -65 -342 21 -319
rect 176 -342 229 -319
rect 646 -320 1045 -319
rect 384 -322 1045 -320
rect 384 -339 690 -322
rect 707 -339 770 -322
rect 787 -339 814 -322
rect 831 -339 898 -322
rect 915 -339 978 -322
rect 995 -339 1022 -322
rect 1039 -339 1045 -322
rect 384 -342 1045 -339
use invx  invx_0
timestamp 1726352782
transform 1 0 117 0 1 -287
box -96 -55 59 239
use invx  invx_1
timestamp 1726352782
transform 1 0 325 0 1 -287
box -96 -55 59 239
use invx  invx_2
timestamp 1726352782
transform 1 0 -89 0 1 58
box -96 -55 59 239
use invx  invx_3
timestamp 1726352782
transform 1 0 -124 0 1 -287
box -96 -55 59 239
use invx  invx_4
timestamp 1726352782
transform 1 0 531 0 1 -287
box -96 -55 59 239
use just_tg  just_tg_0
timestamp 1726407028
transform 1 0 95 0 1 55
box -95 -55 59 228
use just_tg  just_tg_1
timestamp 1726407028
transform -1 0 213 0 1 55
box -95 -55 59 228
<< labels >>
rlabel metal1 682 -331 682 -331 7 vss
port 3 w
rlabel metal1 682 -59 682 -59 7 vdd
port 2 w
rlabel metal1 890 -331 890 -331 7 vss
port 3 w
rlabel metal1 890 -59 890 -59 7 vdd
port 2 w
rlabel metal1 -220 -331 -220 -331 1 Vss
port 8 n
rlabel metal1 -186 286 -186 286 1 Vdd
port 7 n
rlabel locali -131 114 -131 114 1 D
port 5 n
rlabel locali 861 -241 861 -241 5 Q
port 9 s
rlabel locali -166 -231 -166 -231 7 CLK
port 6 w
<< end >>
